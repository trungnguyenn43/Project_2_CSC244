
module project2_csc244();

endmodule